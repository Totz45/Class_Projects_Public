library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity IFID_reg is 
	port( clk       : in  std_logic;
			rst       : in  std_logic; 
			pc4_in:					IN STD_LOGIC_VECTOR(31 downto 0);
			instrMem_in:  					IN STD_LOGIC_VECTOR(31 downto 0);
			pc4_out: 				OUT STD_LOGIC_VECTOR(31 downto 0);
			instrMem_out: 				OUT STD_LOGIC_VECTOR(31 downto 0));
end entity IFID_reg;

architecture Behavioral of IFID_reg is
begin
    process(clk, rst)
    begin
        if rst = '1' then
            -- When reset is high, clear the stored instruction and PC.
            instrMem_out <= (others => '0');
            pc4_out    <= (others => '0');
        elsif rising_edge(clk) then
            -- On each rising edge the IF/ID register captures the values coming from IF stage.
            instrMem_out <= instrMem_in;
            pc4_out    <= pc4_in;
        end if;
    end process;
end Behavioral;


