-- File Name: WriteUnit.vhd
-- Author: Tate Finley
-- Purpose: write only functionality for the registers.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.RegisterPackage.ALL;

entity WriteUnit is
    Port (Clock : in STD_LOGIC;
			reg_write_sig : in STD_LOGIC;
			reg_write_1 : in STD_LOGIC_VECTOR(4 downto 0);
			reg_data : in STD_LOGIC_VECTOR(31 downto 0);
			all_regs_with_data : inout RegisterArrayType);
end WriteUnit;

architecture Structural of WriteUnit is
    signal reg_enable_sig : STD_LOGIC_VECTOR(31 downto 0);
    signal write_enable_sig: STD_LOGIC_VECTOR(31 downto 0);

    -- Components located inside the write section of the register unit
    component Register_decoder
			port(	S: in STD_LOGIC_VECTOR(4 downto 0);
					Z: out STD_LOGIC_VECTOR(31 downto 0));
	 end component;

    component AND_gate
        Port ( x0 : in STD_LOGIC;
               x1 : in STD_LOGIC;
               Y : out STD_LOGIC);
    end component;

    component reg_unit_registers
        Port ( Clock : in STD_LOGIC;
               C : in STD_LOGIC;
               D : in STD_LOGIC_VECTOR(31 downto 0);
               Q : out STD_LOGIC_VECTOR(31 downto 0));
    end component;

begin
    -- Instantiate decoder
    DUT1: Register_decoder port map (reg_write_1,reg_enable_sig);

    -- Generate AND gates and register instances
    Create_Connections: for i in 0 to 31 generate
        DUT2: AND_gate port map (reg_enable_sig(i), reg_write_sig, write_enable_sig(i));

        DUT3: reg_unit_registers port map (Clock, write_enable_sig(i), reg_data, all_regs_with_data(i));
    end generate;

end Structural;
